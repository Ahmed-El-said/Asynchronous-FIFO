module FIFO (
    
);
    
endmodule